hello world pretend this is code

 goodbye world

hello world pretend this is code
